`timescale 1ns/1ps
// 32 bit inputs, 32 bit outputs, ignore overflow, asynchronous
module adder (

);



endmodule