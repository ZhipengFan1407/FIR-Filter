`timescale 1ns/1ps

module distr_arith (
    input clk3
);

endmodule