`timescale 1ns/1ps
// A counter that starts counting from an activation of a signal, and sends out
// an enable signal to the output DFF
module counter(

);



endmodule