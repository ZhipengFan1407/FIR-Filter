`timescale 1ns/1ps
// 32 bit input, 32 bit output, left shift by 1 bit, asynchronous
module left_shift_1(

);



endmodule