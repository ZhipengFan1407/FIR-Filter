`timescale 1ns/1ps
// 32 bit input, 32 bit output, D Flip Flop with Enable feature, Enable is not used for
// the scale accumulation, but the output sum since only output after all 16 bits of
// all inputs are processed
module dff_en(

);



endmodule